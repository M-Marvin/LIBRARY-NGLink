voltage divider netlist
V1 in 0 10
R1 in out 1k
R2 out 0 2k
.end
